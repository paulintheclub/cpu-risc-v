@00000000
93010000 6F000005 23A08101 23A29101 
23A4A101 23A6B101 23A8C101 23AAD101 
23ACE101 23AEF101 93810102 67800000 
130C0000 930C0000 130D0000 930D0000 
130E0000 930E0000 130F0000 930F0000 
67800000 13050010 93050001 131C7501 
93DC8500 135DFC41 930DF5FF 134E0D80 
937E0D80 13EF0D80 971F0000 EFF0DFF8 
13058000 370C8000 13000000 B31CAC00 
335DAC00 B3DDAC40 330EAC00 B3CEBC01 
33FFBC01 B3EFDC01 EFF01FF6 13051000 
9305F0FF 132CF5FF 933CF5FF 33ADA500 
B3BDA500 330EB540 B38EB540 330FA040 
B38FA540 EFF05FF3 13051000 9305000C 
338CA500 B30CAC00 338D8C41 B30DAC41 
23A0BD01 03AE0D00 930ECEFF 03AF4E00 
2322EF01 83AF8E00 EFF01FF0 13052000 
9315E501 338CA502 B3BCA502 339DA502 
B32DAD02 130E000F 939D4D00 93DD4D00 
B32EBE03 338FAE00 B30FEF03 EFF0DFEC 
13050000 9305F0FF 6304B500 930CB007 
6314B500 130DB007 6344B500 930DB007 
6364B500 130EB007 63D4A500 930EB007 
63F4A500 130FB007 EFF01FE9 73001000 
