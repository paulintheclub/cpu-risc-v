@00000000
80000000
00000000
FFFFFFFF
000000FF
000007FF
FFFFF800   
FFFFF8FF
00001078
00800000
80000000
00008000
FF800000
00800008
7F800000
80000000   
FF800000
00000000
00000001
00000001
00000000
00000002
00000000
FFFFFFFF
FFFFFFFE
000000C1
000000C2
00000001
000000C0
000000C0
000000BC
000000C0
000000C0
00000000
00000001
FFFFFFFF
0FFFFFFF
000000F0
0000000E
00000010
00000100
00000000
0000007B
FFFFFFFF
0000007B
000000F0
0000007B
00000010
00000100
000000C0
000000C0
